
module xor_block(input in1,in2,
                     output out1);

assign out1 = in1 ^ in2;

endmodule
